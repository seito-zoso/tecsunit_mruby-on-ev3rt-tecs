import("EV3_common.cdl");
import("TECSInfo.cdl");
//[domain(HRP2, "trusted")]
//[domain(HRP2, "nontrusted")]
celltype tTaskMain {
	entry sTaskBody eBody;

	call sKernel 	cKernel;
	call sLCD 		cLCD;
	call sButton	cButton;

	/* TECSInfo */
  call  nTECSInfo::sTECSInfo cTECSInfo;
  [dynamic,optional]
      call  nTECSInfo::sNamespaceInfo cNSInfo;
  [dynamic,optional]
      call  nTECSInfo::sRegionInfo    cRegionInfo;
  [dynamic,optional]
      call  nTECSInfo::sCellInfo      cCellInfo;
  [dynamic,optional]
      call  nTECSInfo::sSignatureInfo cSignatureInfo;
  [dynamic,optional]
      call  nTECSInfo::sCelltypeInfo  cCelltypeInfo;
  [dynamic,optional]
      call  nTECSInfo::sVarDeclInfo   cVarDeclInfo;
  [dynamic,optional]
      call  nTECSInfo::sTypeInfo      cTypeInfo;
  [dynamic,optional]
      call  nTECSInfo::sFunctionInfo  cFunctionInfo;
  [dynamic,optional]
      call  nTECSInfo::sParamInfo     cParamInfo;
  [dynamic,optional]
      call  nTECSInfo::sEntryInfo     cEntryInfo;

};

region rDomainEV3 {

	cell tTaskMain TaskMain {
		cTECSinfo = TECSInfo.eTECSInfo;

    cKernel = HRP2Kernel.eKernel;
    cButton = Button.eButton;
    cLCD = LCD.eLCD;
	};

	cell tTask Task {
	// 呼び口の結合
		cBody = TaskMain.eBody;
		//* 属性の設定
		taskAttribute 	= C_EXP("TA_ACT");
		priority 		= C_EXP("EV3_MRUBY_VM_PRIORITY");
		systemStackSize = C_EXP("MRUBY_VM_STACK_SIZE");
		//userStackSize = C_EXP("STACK_SIZE");
	};

};
